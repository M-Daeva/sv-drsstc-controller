`include "modules/defines.sv"
`include "modules/pwm.sv"
`include "modules/edge_det.sv"
`include "modules/sync.sv"
