/*
calculates bus width from its max value
`width(255) -> 8
*/
`define width(val) $clog2(val+1)


`define reg(val) reg[$clog2(val+1)-1:0]

`define wire(val) wire[$clog2(val+1)-1:0]

/*
defines 2d array reg
`reg_2d(my_array, 255, 4) -> reg[8] my_array [4:0]
*/
`define reg_2d(name, width_val, length_val) reg[$clog2(width_val+1)-1:0] \
 ``name`` [length_val:0]

/*
defines 2d array wire
`wire_2d(my_array, 255, 4) -> wire[8] my_array [4:0]
*/
`define wire_2d(name, width_val, length_val) wire[$clog2(width_val+1)-1:0] \
 ``name`` [length_val:0]

`define div(A, B) A / B + (2*(A % B) >= B ? 1 : 0)

`define lookup \
8'd1: cnt <= 17'd99999; \
8'd2: cnt <= 17'd49999; \
8'd3: cnt <= 17'd33332; \
8'd4: cnt <= 17'd24999; \
8'd5: cnt <= 17'd19999; \
8'd6: cnt <= 17'd16666; \
8'd7: cnt <= 17'd14285; \
8'd8: cnt <= 17'd12499; \
8'd9: cnt <= 17'd11110; \
8'd10: cnt <= 17'd9999; \
8'd11: cnt <= 17'd9090; \
8'd12: cnt <= 17'd8332; \
8'd13: cnt <= 17'd7691; \
8'd14: cnt <= 17'd7142; \
8'd15: cnt <= 17'd6666; \
8'd16: cnt <= 17'd6249; \
8'd17: cnt <= 17'd5881; \
8'd18: cnt <= 17'd5555; \
8'd19: cnt <= 17'd5262; \
8'd20: cnt <= 17'd4999; \
8'd21: cnt <= 17'd4761; \
8'd22: cnt <= 17'd4544; \
8'd23: cnt <= 17'd4347; \
8'd24: cnt <= 17'd4166; \
8'd25: cnt <= 17'd3999; \
8'd26: cnt <= 17'd3845; \
8'd27: cnt <= 17'd3703; \
8'd28: cnt <= 17'd3570; \
8'd29: cnt <= 17'd3447; \
8'd30: cnt <= 17'd3332; \
8'd31: cnt <= 17'd3225; \
8'd32: cnt <= 17'd3124; \
8'd33: cnt <= 17'd3029; \
8'd34: cnt <= 17'd2940; \
8'd35: cnt <= 17'd2856; \
8'd36: cnt <= 17'd2777; \
8'd37: cnt <= 17'd2702; \
8'd38: cnt <= 17'd2631; \
8'd39: cnt <= 17'd2563; \
8'd40: cnt <= 17'd2499; \
8'd41: cnt <= 17'd2438; \
8'd42: cnt <= 17'd2380; \
8'd43: cnt <= 17'd2325; \
8'd44: cnt <= 17'd2272; \
8'd45: cnt <= 17'd2221; \
8'd46: cnt <= 17'd2173; \
8'd47: cnt <= 17'd2127; \
8'd48: cnt <= 17'd2082; \
8'd49: cnt <= 17'd2040; \
8'd50: cnt <= 17'd1999; \
8'd51: cnt <= 17'd1960; \
8'd52: cnt <= 17'd1922; \
8'd53: cnt <= 17'd1886; \
8'd54: cnt <= 17'd1851; \
8'd55: cnt <= 17'd1817; \
8'd56: cnt <= 17'd1785; \
8'd57: cnt <= 17'd1753; \
8'd58: cnt <= 17'd1723; \
8'd59: cnt <= 17'd1694; \
8'd60: cnt <= 17'd1666; \
8'd61: cnt <= 17'd1638; \
8'd62: cnt <= 17'd1612; \
8'd63: cnt <= 17'd1586; \
8'd64: cnt <= 17'd1562; \
8'd65: cnt <= 17'd1537; \
8'd66: cnt <= 17'd1514; \
8'd67: cnt <= 17'd1492; \
8'd68: cnt <= 17'd1470; \
8'd69: cnt <= 17'd1448; \
8'd70: cnt <= 17'd1428; \
8'd71: cnt <= 17'd1407; \
8'd72: cnt <= 17'd1388; \
8'd73: cnt <= 17'd1369; \
8'd74: cnt <= 17'd1350; \
8'd75: cnt <= 17'd1332; \
8'd76: cnt <= 17'd1315; \
8'd77: cnt <= 17'd1298; \
8'd78: cnt <= 17'd1281; \
8'd79: cnt <= 17'd1265; \
8'd80: cnt <= 17'd1249; \
8'd81: cnt <= 17'd1234; \
8'd82: cnt <= 17'd1219; \
8'd83: cnt <= 17'd1204; \
8'd84: cnt <= 17'd1189; \
8'd85: cnt <= 17'd1175; \
8'd86: cnt <= 17'd1162; \
8'd87: cnt <= 17'd1148; \
8'd88: cnt <= 17'd1135; \
8'd89: cnt <= 17'd1123; \
8'd90: cnt <= 17'd1110; \
8'd91: cnt <= 17'd1098; \
8'd92: cnt <= 17'd1086; \
8'd93: cnt <= 17'd1074; \
8'd94: cnt <= 17'd1063; \
8'd95: cnt <= 17'd1052; \
8'd96: cnt <= 17'd1041; \
8'd97: cnt <= 17'd1030; \
8'd98: cnt <= 17'd1019; \
8'd99: cnt <= 17'd1009; \
8'd100: cnt <= 17'd999; \
8'd101: cnt <= 17'd989; \
8'd102: cnt <= 17'd979; \
8'd103: cnt <= 17'd970; \
8'd104: cnt <= 17'd961; \
8'd105: cnt <= 17'd951; \
8'd106: cnt <= 17'd942; \
8'd107: cnt <= 17'd934; \
8'd108: cnt <= 17'd925; \
8'd109: cnt <= 17'd916; \
8'd110: cnt <= 17'd908; \
8'd111: cnt <= 17'd900; \
8'd112: cnt <= 17'd892; \
8'd113: cnt <= 17'd884; \
8'd114: cnt <= 17'd876; \
8'd115: cnt <= 17'd869; \
8'd116: cnt <= 17'd861; \
8'd117: cnt <= 17'd854; \
8'd118: cnt <= 17'd846; \
8'd119: cnt <= 17'd839; \
8'd120: cnt <= 17'd832; \
8'd121: cnt <= 17'd825; \
8'd122: cnt <= 17'd819; \
8'd123: cnt <= 17'd812; \
8'd124: cnt <= 17'd805; \
8'd125: cnt <= 17'd799; \
8'd126: cnt <= 17'd793; \
8'd127: cnt <= 17'd786; \
8'd128: cnt <= 17'd780; \
8'd129: cnt <= 17'd774; \
8'd130: cnt <= 17'd768; \
8'd131: cnt <= 17'd762; \
8'd132: cnt <= 17'd757; \
8'd133: cnt <= 17'd751; \
8'd134: cnt <= 17'd745; \
8'd135: cnt <= 17'd740; \
8'd136: cnt <= 17'd734; \
8'd137: cnt <= 17'd729; \
8'd138: cnt <= 17'd724; \
8'd139: cnt <= 17'd718; \
8'd140: cnt <= 17'd713; \
8'd141: cnt <= 17'd708; \
8'd142: cnt <= 17'd703; \
8'd143: cnt <= 17'd698; \
8'd144: cnt <= 17'd693; \
8'd145: cnt <= 17'd689; \
8'd146: cnt <= 17'd684; \
8'd147: cnt <= 17'd679; \
8'd148: cnt <= 17'd675; \
8'd149: cnt <= 17'd670; \
8'd150: cnt <= 17'd666; \
8'd151: cnt <= 17'd661; \
8'd152: cnt <= 17'd657; \
8'd153: cnt <= 17'd653; \
8'd154: cnt <= 17'd648; \
8'd155: cnt <= 17'd644; \
8'd156: cnt <= 17'd640; \
8'd157: cnt <= 17'd636; \
8'd158: cnt <= 17'd632; \
8'd159: cnt <= 17'd628; \
8'd160: cnt <= 17'd624; \
8'd161: cnt <= 17'd620; \
8'd162: cnt <= 17'd616; \
8'd163: cnt <= 17'd612; \
8'd164: cnt <= 17'd609; \
8'd165: cnt <= 17'd605; \
8'd166: cnt <= 17'd601; \
8'd167: cnt <= 17'd598; \
8'd168: cnt <= 17'd594; \
8'd169: cnt <= 17'd591; \
8'd170: cnt <= 17'd587; \
8'd171: cnt <= 17'd584; \
8'd172: cnt <= 17'd580; \
8'd173: cnt <= 17'd577; \
8'd174: cnt <= 17'd574; \
8'd175: cnt <= 17'd570; \
8'd176: cnt <= 17'd567; \
8'd177: cnt <= 17'd564; \
8'd178: cnt <= 17'd561; \
8'd179: cnt <= 17'd558; \
8'd180: cnt <= 17'd555; \
8'd181: cnt <= 17'd551; \
8'd182: cnt <= 17'd548; \
8'd183: cnt <= 17'd545; \
8'd184: cnt <= 17'd542; \
8'd185: cnt <= 17'd540; \
8'd186: cnt <= 17'd537; \
8'd187: cnt <= 17'd534; \
8'd188: cnt <= 17'd531; \
8'd189: cnt <= 17'd528; \
8'd190: cnt <= 17'd525; \
8'd191: cnt <= 17'd523; \
8'd192: cnt <= 17'd520; \
8'd193: cnt <= 17'd517; \
8'd194: cnt <= 17'd514; \
8'd195: cnt <= 17'd512; \
8'd196: cnt <= 17'd509; \
8'd197: cnt <= 17'd507; \
8'd198: cnt <= 17'd504; \
8'd199: cnt <= 17'd502; \
8'd200: cnt <= 17'd499; \
8'd201: cnt <= 17'd497; \
8'd202: cnt <= 17'd494; \
8'd203: cnt <= 17'd492; \
8'd204: cnt <= 17'd489; \
8'd205: cnt <= 17'd487; \
8'd206: cnt <= 17'd484; \
8'd207: cnt <= 17'd482; \
8'd208: cnt <= 17'd480; \
8'd209: cnt <= 17'd477; \
8'd210: cnt <= 17'd475; \
8'd211: cnt <= 17'd473; \
8'd212: cnt <= 17'd471; \
8'd213: cnt <= 17'd468; \
8'd214: cnt <= 17'd466; \
8'd215: cnt <= 17'd464; \
8'd216: cnt <= 17'd462; \
8'd217: cnt <= 17'd460; \
8'd218: cnt <= 17'd458; \
8'd219: cnt <= 17'd456; \
8'd220: cnt <= 17'd454; \
8'd221: cnt <= 17'd451; \
8'd222: cnt <= 17'd449; \
8'd223: cnt <= 17'd447; \
8'd224: cnt <= 17'd445; \
8'd225: cnt <= 17'd443; \
8'd226: cnt <= 17'd441; \
8'd227: cnt <= 17'd440; \
8'd228: cnt <= 17'd438; \
8'd229: cnt <= 17'd436; \
8'd230: cnt <= 17'd434; \
8'd231: cnt <= 17'd432; \
8'd232: cnt <= 17'd430; \
8'd233: cnt <= 17'd428; \
8'd234: cnt <= 17'd426; \
8'd235: cnt <= 17'd425; \
8'd236: cnt <= 17'd423; \
8'd237: cnt <= 17'd421; \
8'd238: cnt <= 17'd419; \
8'd239: cnt <= 17'd417; \
8'd240: cnt <= 17'd416; \
8'd241: cnt <= 17'd414; \
8'd242: cnt <= 17'd412; \
8'd243: cnt <= 17'd411; \
8'd244: cnt <= 17'd409; \
8'd245: cnt <= 17'd407; \
8'd246: cnt <= 17'd406; \
8'd247: cnt <= 17'd404; \
8'd248: cnt <= 17'd402; \
8'd249: cnt <= 17'd401; \
8'd250: cnt <= 17'd399; \
8'd251: cnt <= 17'd397; \
8'd252: cnt <= 17'd396; \
8'd253: cnt <= 17'd394; \
8'd254: cnt <= 17'd393; \
8'd255: cnt <= 17'd391;
