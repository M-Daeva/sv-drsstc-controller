/*
calculates bus width from its max value
`width(255) -> 8
*/
`define width(val) $clog2(val+1)


`define reg(val) reg[$clog2(val+1)-1:0]

`define wire(val) wire[$clog2(val+1)-1:0]

/*
defines 2d array reg
`reg_2d(my_array, 255, 4) -> reg[8] my_array [4:0]
*/
`define reg_2d(name, width_val, length_val) reg[$clog2(width_val+1)-1:0] \
 ``name`` [length_val:0]

/*
defines 2d array wire
`wire_2d(my_array, 255, 4) -> wire[8] my_array [4:0]
*/
`define wire_2d(name, width_val, length_val) wire[$clog2(width_val+1)-1:0] \
 ``name`` [length_val:0]

`define div(A, B) A / B + (2*(A % B) >= B ? 1 : 0)

`define lookup \
8'd1: cnt <= 14'd9999; \
8'd2: cnt <= 14'd4999; \
8'd3: cnt <= 14'd3332; \
8'd4: cnt <= 14'd2499; \
8'd5: cnt <= 14'd1999; \
8'd6: cnt <= 14'd1666; \
8'd7: cnt <= 14'd1428; \
8'd8: cnt <= 14'd1249; \
8'd9: cnt <= 14'd1110; \
8'd10: cnt <= 14'd999; \
8'd11: cnt <= 14'd908; \
8'd12: cnt <= 14'd832; \
8'd13: cnt <= 14'd768; \
8'd14: cnt <= 14'd713; \
8'd15: cnt <= 14'd666; \
8'd16: cnt <= 14'd624; \
8'd17: cnt <= 14'd587; \
8'd18: cnt <= 14'd555; \
8'd19: cnt <= 14'd525; \
8'd20: cnt <= 14'd499; \
8'd21: cnt <= 14'd475; \
8'd22: cnt <= 14'd454; \
8'd23: cnt <= 14'd434; \
8'd24: cnt <= 14'd416; \
8'd25: cnt <= 14'd399; \
8'd26: cnt <= 14'd384; \
8'd27: cnt <= 14'd369; \
8'd28: cnt <= 14'd356; \
8'd29: cnt <= 14'd344; \
8'd30: cnt <= 14'd332; \
8'd31: cnt <= 14'd322; \
8'd32: cnt <= 14'd312; \
8'd33: cnt <= 14'd302; \
8'd34: cnt <= 14'd293; \
8'd35: cnt <= 14'd285; \
8'd36: cnt <= 14'd277; \
8'd37: cnt <= 14'd269; \
8'd38: cnt <= 14'd262; \
8'd39: cnt <= 14'd255; \
8'd40: cnt <= 14'd249; \
8'd41: cnt <= 14'd243; \
8'd42: cnt <= 14'd237; \
8'd43: cnt <= 14'd232; \
8'd44: cnt <= 14'd226; \
8'd45: cnt <= 14'd221; \
8'd46: cnt <= 14'd216; \
8'd47: cnt <= 14'd212; \
8'd48: cnt <= 14'd207; \
8'd49: cnt <= 14'd203; \
8'd50: cnt <= 14'd199; \
8'd51: cnt <= 14'd195; \
8'd52: cnt <= 14'd191; \
8'd53: cnt <= 14'd188; \
8'd54: cnt <= 14'd184; \
8'd55: cnt <= 14'd181; \
8'd56: cnt <= 14'd178; \
8'd57: cnt <= 14'd174; \
8'd58: cnt <= 14'd171; \
8'd59: cnt <= 14'd168; \
8'd60: cnt <= 14'd166; \
8'd61: cnt <= 14'd163; \
8'd62: cnt <= 14'd160; \
8'd63: cnt <= 14'd158; \
8'd64: cnt <= 14'd155; \
8'd65: cnt <= 14'd153; \
8'd66: cnt <= 14'd151; \
8'd67: cnt <= 14'd148; \
8'd68: cnt <= 14'd146; \
8'd69: cnt <= 14'd144; \
8'd70: cnt <= 14'd142; \
8'd71: cnt <= 14'd140; \
8'd72: cnt <= 14'd138; \
8'd73: cnt <= 14'd136; \
8'd74: cnt <= 14'd134; \
8'd75: cnt <= 14'd132; \
8'd76: cnt <= 14'd131; \
8'd77: cnt <= 14'd129; \
8'd78: cnt <= 14'd127; \
8'd79: cnt <= 14'd126; \
8'd80: cnt <= 14'd124; \
8'd81: cnt <= 14'd122; \
8'd82: cnt <= 14'd121; \
8'd83: cnt <= 14'd119; \
8'd84: cnt <= 14'd118; \
8'd85: cnt <= 14'd117; \
8'd86: cnt <= 14'd115; \
8'd87: cnt <= 14'd114; \
8'd88: cnt <= 14'd113; \
8'd89: cnt <= 14'd111; \
8'd90: cnt <= 14'd110; \
8'd91: cnt <= 14'd109; \
8'd92: cnt <= 14'd108; \
8'd93: cnt <= 14'd107; \
8'd94: cnt <= 14'd105; \
8'd95: cnt <= 14'd104; \
8'd96: cnt <= 14'd103; \
8'd97: cnt <= 14'd102; \
8'd98: cnt <= 14'd101; \
8'd99: cnt <= 14'd100; \
8'd100: cnt <= 14'd99; \
8'd101: cnt <= 14'd98; \
8'd102: cnt <= 14'd97; \
8'd103: cnt <= 14'd96; \
8'd104: cnt <= 14'd95; \
8'd105: cnt <= 14'd94; \
8'd106: cnt <= 14'd93; \
8'd107: cnt <= 14'd92; \
8'd108: cnt <= 14'd92; \
8'd109: cnt <= 14'd91; \
8'd110: cnt <= 14'd90; \
8'd111: cnt <= 14'd89; \
8'd112: cnt <= 14'd88; \
8'd113: cnt <= 14'd87; \
8'd114: cnt <= 14'd87; \
8'd115: cnt <= 14'd86; \
8'd116: cnt <= 14'd85; \
8'd117: cnt <= 14'd84; \
8'd118: cnt <= 14'd84; \
8'd119: cnt <= 14'd83; \
8'd120: cnt <= 14'd82; \
8'd121: cnt <= 14'd82; \
8'd122: cnt <= 14'd81; \
8'd123: cnt <= 14'd80; \
8'd124: cnt <= 14'd80; \
8'd125: cnt <= 14'd79; \
8'd126: cnt <= 14'd78; \
8'd127: cnt <= 14'd78; \
8'd128: cnt <= 14'd77; \
8'd129: cnt <= 14'd77; \
8'd130: cnt <= 14'd76; \
8'd131: cnt <= 14'd75; \
8'd132: cnt <= 14'd75; \
8'd133: cnt <= 14'd74; \
8'd134: cnt <= 14'd74; \
8'd135: cnt <= 14'd73; \
8'd136: cnt <= 14'd73; \
8'd137: cnt <= 14'd72; \
8'd138: cnt <= 14'd71; \
8'd139: cnt <= 14'd71; \
8'd140: cnt <= 14'd70; \
8'd141: cnt <= 14'd70; \
8'd142: cnt <= 14'd69; \
8'd143: cnt <= 14'd69; \
8'd144: cnt <= 14'd68; \
8'd145: cnt <= 14'd68; \
8'd146: cnt <= 14'd67; \
8'd147: cnt <= 14'd67; \
8'd148: cnt <= 14'd67; \
8'd149: cnt <= 14'd66; \
8'd150: cnt <= 14'd66; \
8'd151: cnt <= 14'd65; \
8'd152: cnt <= 14'd65; \
8'd153: cnt <= 14'd64; \
8'd154: cnt <= 14'd64; \
8'd155: cnt <= 14'd64; \
8'd156: cnt <= 14'd63; \
8'd157: cnt <= 14'd63; \
8'd158: cnt <= 14'd62; \
8'd159: cnt <= 14'd62; \
8'd160: cnt <= 14'd62; \
8'd161: cnt <= 14'd61; \
8'd162: cnt <= 14'd61; \
8'd163: cnt <= 14'd60; \
8'd164: cnt <= 14'd60; \
8'd165: cnt <= 14'd60; \
8'd166: cnt <= 14'd59; \
8'd167: cnt <= 14'd59; \
8'd168: cnt <= 14'd59; \
8'd169: cnt <= 14'd58; \
8'd170: cnt <= 14'd58; \
8'd171: cnt <= 14'd57; \
8'd172: cnt <= 14'd57; \
8'd173: cnt <= 14'd57; \
8'd174: cnt <= 14'd56; \
8'd175: cnt <= 14'd56; \
8'd176: cnt <= 14'd56; \
8'd177: cnt <= 14'd55; \
8'd178: cnt <= 14'd55; \
8'd179: cnt <= 14'd55; \
8'd180: cnt <= 14'd55; \
8'd181: cnt <= 14'd54; \
8'd182: cnt <= 14'd54; \
8'd183: cnt <= 14'd54; \
8'd184: cnt <= 14'd53; \
8'd185: cnt <= 14'd53; \
8'd186: cnt <= 14'd53; \
8'd187: cnt <= 14'd52; \
8'd188: cnt <= 14'd52; \
8'd189: cnt <= 14'd52; \
8'd190: cnt <= 14'd52; \
8'd191: cnt <= 14'd51; \
8'd192: cnt <= 14'd51; \
8'd193: cnt <= 14'd51; \
8'd194: cnt <= 14'd51; \
8'd195: cnt <= 14'd50; \
8'd196: cnt <= 14'd50; \
8'd197: cnt <= 14'd50; \
8'd198: cnt <= 14'd50; \
8'd199: cnt <= 14'd49; \
8'd200: cnt <= 14'd49; \
8'd201: cnt <= 14'd49; \
8'd202: cnt <= 14'd49; \
8'd203: cnt <= 14'd48; \
8'd204: cnt <= 14'd48; \
8'd205: cnt <= 14'd48; \
8'd206: cnt <= 14'd48; \
8'd207: cnt <= 14'd47; \
8'd208: cnt <= 14'd47; \
8'd209: cnt <= 14'd47; \
8'd210: cnt <= 14'd47; \
8'd211: cnt <= 14'd46; \
8'd212: cnt <= 14'd46; \
8'd213: cnt <= 14'd46; \
8'd214: cnt <= 14'd46; \
8'd215: cnt <= 14'd46; \
8'd216: cnt <= 14'd45; \
8'd217: cnt <= 14'd45; \
8'd218: cnt <= 14'd45; \
8'd219: cnt <= 14'd45; \
8'd220: cnt <= 14'd44; \
8'd221: cnt <= 14'd44; \
8'd222: cnt <= 14'd44; \
8'd223: cnt <= 14'd44; \
8'd224: cnt <= 14'd44; \
8'd225: cnt <= 14'd43; \
8'd226: cnt <= 14'd43; \
8'd227: cnt <= 14'd43; \
8'd228: cnt <= 14'd43; \
8'd229: cnt <= 14'd43; \
8'd230: cnt <= 14'd42; \
8'd231: cnt <= 14'd42; \
8'd232: cnt <= 14'd42; \
8'd233: cnt <= 14'd42; \
8'd234: cnt <= 14'd42; \
8'd235: cnt <= 14'd42; \
8'd236: cnt <= 14'd41; \
8'd237: cnt <= 14'd41; \
8'd238: cnt <= 14'd41; \
8'd239: cnt <= 14'd41; \
8'd240: cnt <= 14'd41; \
8'd241: cnt <= 14'd40; \
8'd242: cnt <= 14'd40; \
8'd243: cnt <= 14'd40; \
8'd244: cnt <= 14'd40; \
8'd245: cnt <= 14'd40; \
8'd246: cnt <= 14'd40; \
8'd247: cnt <= 14'd39; \
8'd248: cnt <= 14'd39; \
8'd249: cnt <= 14'd39; \
8'd250: cnt <= 14'd39; \
8'd251: cnt <= 14'd39; \
8'd252: cnt <= 14'd39; \
8'd253: cnt <= 14'd39; \
8'd254: cnt <= 14'd38; \
8'd255: cnt <= 14'd38;
